package DummyWriteEnvPkg;
endpackage
