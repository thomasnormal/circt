// Wrapper to inject prim_assert macros for usbdev_aon_wake.
`include "prim_assert.sv"
`include "usbdev_aon_wake.sv"
