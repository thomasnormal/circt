module ovl_sem_next(input logic clk);
  logic reset = 1'b1;
  logic enable = 1'b1;
  logic start_event = 1'b1;
`ifdef FAIL
  logic test_expr = 1'b0;
`else
  logic test_expr = 1'b1;
`endif
  ovl_next #(
      .num_cks(1),
      .check_overlapping(1),
      .check_missing_start(0)) dut (
      .clock(clk),
      .reset(reset),
      .enable(enable),
      .start_event(start_event),
      .test_expr(test_expr),
      .fire());
endmodule
