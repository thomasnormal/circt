package DummySlaveWriteEnvPkg;
endpackage
