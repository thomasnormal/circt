`vendor_directive foo bar baz
module top;
endmodule
