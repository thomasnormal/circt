// RUN: circt-verilog --ir-moore --no-uvm-auto-include %s 2>&1 | FileCheck %s
// REQUIRES: slang

// Test that $changed is lowered to a sequence-compatible value in concatenation.

module PropertyConcatError(input logic clk, a, b);
  wire x = 'x;

  // $changed uses moore.past to track previous value.
  // CHECK: moore.past
  // CHECK: moore.case_eq
  // CHECK: moore.not
  // CHECK: ltl.concat
  assume property (@(posedge clk) b !== x ##1 $changed(b));

endmodule
