`define HELLO
