module test_finish;
  initial begin
    $display("About to finish");
    $finish;
  end
endmodule
