`define WHICH local_cfg_mod
