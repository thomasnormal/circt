// RUN: circt-verilog %s --ir-moore | FileCheck %s

module CrossSelectSetExprFunctionCasePushbackSupported;
  bit clk;
  bit [1:0] a, b;

  covergroup cg @(posedge clk);
    coverpoint a;
    coverpoint b;
    X: cross a, b {
      function CrossQueueType mk(int lim);
        case (lim)
          0: mk.push_back('{0, 0});
          1: mk.push_back('{1, 1});
          default: begin
            mk.push_back('{0, 1});
            mk.push_back('{1, 0});
          end
        endcase
      endfunction
      bins one = mk(2);
    }
  endgroup
endmodule

// CHECK: moore.crossbin.decl @one kind<bins> {
// CHECK:   moore.binsof @a intersect [0]
// CHECK:   moore.binsof @b intersect [1]
// CHECK:   moore.binsof @a intersect [1] {group = 1 : i32}
// CHECK:   moore.binsof @b intersect [0] {group = 1 : i32}
// CHECK: }
