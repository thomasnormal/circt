module top;
  helper u();
endmodule
