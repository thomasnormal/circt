// Wrapper to inject prim_assert macros for usb_fs_nb_out_pe.
`include "prim_assert.sv"
`include "usb_fs_nb_out_pe.sv"
