`include "cfg.svh"
module `WHICH;
endmodule
