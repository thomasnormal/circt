// RUN: circt-verilog --parse-only --no-uvm-auto-include -I ~/uvm-core/src ~/uvm-core/src/uvm_pkg.sv %s
// RUN: circt-verilog --ir-moore --no-uvm-auto-include -I ~/uvm-core/src ~/uvm-core/src/uvm_pkg.sv %s | FileCheck %s --check-prefix=MOORE
// REQUIRES: slang
// XFAIL: *
// Currently trips always_ff driver legality checks in imported UVM code.

//===----------------------------------------------------------------------===//
// AVIP End-to-End Testbench - Iteration 63 Track A
//===----------------------------------------------------------------------===//
//
// This testbench demonstrates a complete AVIP-style verification environment
// using the CIRCT UVM stubs. It exercises:
//
// 1. UVM component hierarchy (env, agent, driver, monitor, sequencer)
// 2. Virtual interface with timing (@posedge clk)
// 3. Randomization with constraints
// 4. Coverage collection with covergroups
// 5. TLM communication (analysis ports)
//
// This represents the target for CIRCT UVM parity with commercial simulators.
//
//===----------------------------------------------------------------------===//
//
// STATUS (Iteration 63):
//   - Parsing: PASS (all UVM components parse correctly)
//   - Moore IR: PASS (all constructs convert to Moore IR)
//   - Full Lowering: BLOCKED (timing in class tasks needs process context)
//
// KNOWN LIMITATIONS:
//   1. Type cast of virtual interface signals not fully supported
//      Workaround: Use if/else with direct enum assignment
//   2. Timing controls (@posedge, #delay) in class tasks require llhd.process
//      This is the main blocker for full LLHD lowering
//   3. Clocking blocks and modports with virtual interfaces have limited support
//      Workaround: Use direct interface signal access
//
// WHAT WORKS:
//   - UVM class hierarchy with inheritance
//   - Virtual interface access in class methods
//   - Randomization with constraints (rand, constraint blocks)
//   - Covergroups with coverpoints and cross coverage
//   - Analysis ports and TLM connections
//   - Factory pattern with type_id::create
//   - uvm_config_db access
//
//===----------------------------------------------------------------------===//

`timescale 1ns/1ps
`include "uvm_macros.svh"

//===----------------------------------------------------------------------===//
// Package: APB Protocol Types
//===----------------------------------------------------------------------===//

package avip_apb_pkg;

  // Transfer direction
  typedef enum bit {
    APB_READ  = 1'b0,
    APB_WRITE = 1'b1
  } apb_dir_e;

  // Response status
  typedef enum bit {
    APB_OKAY  = 1'b0,
    APB_ERROR = 1'b1
  } apb_resp_e;

  // Configuration parameters
  parameter int APB_ADDR_W = 32;
  parameter int APB_DATA_W = 32;
  parameter int APB_STRB_W = APB_DATA_W / 8;

endpackage : avip_apb_pkg

// PARSE: module {
// MOORE: module {

//===----------------------------------------------------------------------===//
// Interface: APB Bus Interface
//===----------------------------------------------------------------------===//

interface apb_if (input bit clk, input bit rst_n);
  import avip_apb_pkg::*;

  // APB signals (using bit instead of logic for better virtual interface support)
  bit [APB_ADDR_W-1:0] paddr;
  bit                  pselx;
  bit                  penable;
  bit                  pwrite;
  bit [APB_DATA_W-1:0] pwdata;
  bit [APB_STRB_W-1:0] pstrb;
  bit [APB_DATA_W-1:0] prdata;
  bit                  pready;
  bit                  pslverr;

  // Note: Clocking blocks and modports with virtual interfaces have limited
  // support in CIRCT. Using direct signal access for this test.

endinterface : apb_if

// PARSE-DAG: moore.interface @apb_if
// MOORE-DAG: moore.interface @apb_if

//===----------------------------------------------------------------------===//
// Transaction: APB Sequence Item
//===----------------------------------------------------------------------===//

import uvm_pkg::*;
import avip_apb_pkg::*;

class apb_seq_item extends uvm_sequence_item;
  `uvm_object_utils(apb_seq_item)

  // Random stimulus fields
  rand bit [APB_ADDR_W-1:0] addr;
  rand bit [APB_DATA_W-1:0] wdata;
  rand apb_dir_e            dir;
  rand bit [APB_STRB_W-1:0] strb;

  // Response fields (not randomized)
  bit [APB_DATA_W-1:0] rdata;
  apb_resp_e           resp;

  // Transaction metadata
  int unsigned txn_id;
  static int unsigned txn_counter = 0;

  // Constraints
  constraint c_addr_aligned {
    addr[1:0] == 2'b00;  // Word aligned
  }

  constraint c_addr_range {
    addr[31:8] == 24'b0;  // Limited address space
  }

  constraint c_strb_write {
    dir == APB_WRITE -> strb != 0;  // At least one strobe on write
  }

  constraint c_strb_read {
    dir == APB_READ -> strb == 4'b1111;  // Full word read
  }

  // Constructor
  function new(string name = "apb_seq_item");
    super.new(name);
    txn_id = txn_counter++;
  endfunction

  // Convert to string
  virtual function string convert2string();
    return $sformatf("TXN[%0d] %s addr=0x%08h data=0x%08h strb=%04b",
                     txn_id,
                     dir == APB_WRITE ? "WR" : "RD",
                     addr,
                     dir == APB_WRITE ? wdata : rdata,
                     strb);
  endfunction

  // Copy
  virtual function void do_copy(uvm_object rhs);
    apb_seq_item rhs_item;
    super.do_copy(rhs);
    if ($cast(rhs_item, rhs)) begin
      addr   = rhs_item.addr;
      wdata  = rhs_item.wdata;
      dir    = rhs_item.dir;
      strb   = rhs_item.strb;
      rdata  = rhs_item.rdata;
      resp   = rhs_item.resp;
      txn_id = rhs_item.txn_id;
    end
  endfunction

  // Compare
  virtual function bit do_compare(uvm_object rhs, uvm_comparer comparer);
    apb_seq_item rhs_item;
    if (!$cast(rhs_item, rhs)) return 0;
    return (addr == rhs_item.addr) &&
           (dir == rhs_item.dir) &&
           ((dir == APB_WRITE) ? (wdata == rhs_item.wdata) : 1) &&
           (strb == rhs_item.strb);
  endfunction

endclass : apb_seq_item

// PARSE-DAG: moore.class
// MOORE-DAG: moore.class.classdecl @apb_seq_item

//===----------------------------------------------------------------------===//
// Sequence: APB Base Sequence
//===----------------------------------------------------------------------===//

class apb_base_seq extends uvm_sequence #(apb_seq_item);
  `uvm_object_utils(apb_base_seq)

  // Number of transactions to generate
  rand int unsigned num_txns;

  constraint c_num_txns {
    num_txns inside {[1:20]};
  }

  function new(string name = "apb_base_seq");
    super.new(name);
  endfunction

  virtual task body();
    apb_seq_item item;
    for (int i = 0; i < num_txns; i++) begin
      item = apb_seq_item::type_id::create($sformatf("item_%0d", i));
      start_item(item);
      if (!item.randomize()) begin
        `uvm_error("SEQ", "Randomization failed")
      end
      finish_item(item);
      `uvm_info("SEQ", item.convert2string(), UVM_MEDIUM)
    end
  endtask

endclass : apb_base_seq

//===----------------------------------------------------------------------===//
// Sequencer: APB Sequencer
//===----------------------------------------------------------------------===//

class apb_sequencer extends uvm_sequencer #(apb_seq_item);
  `uvm_component_utils(apb_sequencer)

  function new(string name = "apb_sequencer", uvm_component parent = null);
    super.new(name, parent);
  endfunction

endclass : apb_sequencer

//===----------------------------------------------------------------------===//
// Driver: APB Driver
//===----------------------------------------------------------------------===//

class apb_driver extends uvm_driver #(apb_seq_item);
  `uvm_component_utils(apb_driver)

  // Virtual interface handle (using full interface, not modport)
  virtual apb_if vif;

  function new(string name = "apb_driver", uvm_component parent = null);
    super.new(name, parent);
  endfunction

  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    if (!uvm_config_db#(virtual apb_if)::get(this, "", "vif", vif)) begin
      `uvm_fatal("DRV", "Failed to get virtual interface")
    end
  endfunction

  virtual task run_phase(uvm_phase phase);
    apb_seq_item item;

    // Wait for reset
    @(posedge vif.rst_n);
    `uvm_info("DRV", "Reset released, starting driver", UVM_MEDIUM)

    forever begin
      // Get next item from sequencer
      seq_item_port.get_next_item(req);
      `uvm_info("DRV", {"Driving: ", req.convert2string()}, UVM_HIGH)

      // Drive SETUP phase
      @(posedge vif.clk);
      vif.paddr   <= req.addr;
      vif.pselx   <= 1'b1;
      vif.penable <= 1'b0;
      vif.pwrite  <= (req.dir == APB_WRITE);
      if (req.dir == APB_WRITE) begin
        vif.pwdata <= req.wdata;
        vif.pstrb  <= req.strb;
      end

      // Drive ACCESS phase
      @(posedge vif.clk);
      vif.penable <= 1'b1;

      // Wait for pready
      while (!vif.pready) begin
        @(posedge vif.clk);
      end

      // Capture response
      if (req.dir == APB_READ) begin
        req.rdata = vif.prdata;
      end
      // Note: Type cast of virtual interface signal not fully supported yet
      // Using direct assignment with implicit conversion
      if (vif.pslverr)
        req.resp = APB_ERROR;
      else
        req.resp = APB_OKAY;

      // Return to IDLE
      @(posedge vif.clk);
      vif.pselx   <= 1'b0;
      vif.penable <= 1'b0;

      seq_item_port.item_done();
    end
  endtask

endclass : apb_driver

//===----------------------------------------------------------------------===//
// Monitor: APB Monitor
//===----------------------------------------------------------------------===//

class apb_monitor extends uvm_monitor;
  `uvm_component_utils(apb_monitor)

  // Virtual interface handle (using full interface, not modport)
  virtual apb_if vif;

  // Analysis port for observed transactions
  uvm_analysis_port #(apb_seq_item) analysis_port;

  function new(string name = "apb_monitor", uvm_component parent = null);
    super.new(name, parent);
    analysis_port = new("analysis_port", this);
  endfunction

  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    if (!uvm_config_db#(virtual apb_if)::get(this, "", "vif", vif)) begin
      `uvm_fatal("MON", "Failed to get virtual interface")
    end
  endfunction

  virtual task run_phase(uvm_phase phase);
    apb_seq_item item;

    // Wait for reset
    @(posedge vif.rst_n);
    `uvm_info("MON", "Reset released, starting monitor", UVM_MEDIUM)

    forever begin
      // Wait for valid transaction (psel && penable && pready)
      @(posedge vif.clk);
      if (vif.pselx && vif.penable && vif.pready) begin
        item = apb_seq_item::type_id::create("mon_item");
        item.addr  = vif.paddr;
        // Note: Type cast of virtual interface signal not fully supported
        if (vif.pwrite)
          item.dir = APB_WRITE;
        else
          item.dir = APB_READ;
        item.strb  = vif.pstrb;
        if (item.dir == APB_WRITE) begin
          item.wdata = vif.pwdata;
        end else begin
          item.rdata = vif.prdata;
        end
        // Note: Type cast of virtual interface signal not fully supported
        if (vif.pslverr)
          item.resp = APB_ERROR;
        else
          item.resp = APB_OKAY;

        `uvm_info("MON", {"Observed: ", item.convert2string()}, UVM_HIGH)
        analysis_port.write(item);
      end
    end
  endtask

endclass : apb_monitor

//===----------------------------------------------------------------------===//
// Coverage: APB Functional Coverage
//===----------------------------------------------------------------------===//

class apb_coverage extends uvm_subscriber #(apb_seq_item);
  `uvm_component_utils(apb_coverage)

  // Coverage variables
  bit [APB_ADDR_W-1:0] cov_addr;
  apb_dir_e            cov_dir;
  bit [APB_STRB_W-1:0] cov_strb;
  apb_resp_e           cov_resp;

  // Covergroup
  covergroup apb_cg;
    cp_addr: coverpoint cov_addr[7:2] {
      bins low_addr[]  = {[0:15]};
      bins high_addr[] = {[16:63]};
    }

    cp_dir: coverpoint cov_dir {
      bins read  = {APB_READ};
      bins write = {APB_WRITE};
    }

    cp_strb: coverpoint cov_strb {
      bins full_word   = {4'b1111};
      bins half_word[] = {4'b0011, 4'b1100};
      bins byte_en[]   = {4'b0001, 4'b0010, 4'b0100, 4'b1000};
    }

    cp_resp: coverpoint cov_resp {
      bins okay  = {APB_OKAY};
      bins error = {APB_ERROR};
    }

    // Cross coverage
    addr_x_dir: cross cp_addr, cp_dir;
    dir_x_strb: cross cp_dir, cp_strb {
      ignore_bins read_strb = binsof(cp_dir.read);
    }
  endgroup

  function new(string name = "apb_coverage", uvm_component parent = null);
    super.new(name, parent);
    apb_cg = new();
  endfunction

  // Receive transaction from analysis port
  virtual function void write(apb_seq_item t);
    cov_addr = t.addr;
    cov_dir  = t.dir;
    cov_strb = t.strb;
    cov_resp = t.resp;
    apb_cg.sample();
    `uvm_info("COV", $sformatf("Sampled coverage for %s", t.convert2string()), UVM_HIGH)
  endfunction

  function void report_phase(uvm_phase phase);
    super.report_phase(phase);
    `uvm_info("COV", "Coverage collection complete", UVM_LOW)
  endfunction

endclass : apb_coverage

//===----------------------------------------------------------------------===//
// Agent: APB Agent (Active/Passive)
//===----------------------------------------------------------------------===//

class apb_agent extends uvm_agent;
  `uvm_component_utils(apb_agent)

  // Sub-components
  apb_sequencer sequencer;
  apb_driver    driver;
  apb_monitor   monitor;
  apb_coverage  coverage;

  // Configuration
  bit is_active = 1;

  function new(string name = "apb_agent", uvm_component parent = null);
    super.new(name, parent);
  endfunction

  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);

    // Always build monitor and coverage
    monitor  = apb_monitor::type_id::create("monitor", this);
    coverage = apb_coverage::type_id::create("coverage", this);

    // Build driver and sequencer for active agent
    if (is_active) begin
      sequencer = apb_sequencer::type_id::create("sequencer", this);
      driver    = apb_driver::type_id::create("driver", this);
    end
  endfunction

  virtual function void connect_phase(uvm_phase phase);
    super.connect_phase(phase);

    // Connect monitor to coverage
    monitor.analysis_port.connect(coverage.analysis_export);

    // Connect driver to sequencer for active agent
    if (is_active) begin
      driver.seq_item_port.connect(sequencer.seq_item_export);
    end
  endfunction

endclass : apb_agent

//===----------------------------------------------------------------------===//
// Scoreboard: APB Scoreboard
//===----------------------------------------------------------------------===//

class apb_scoreboard extends uvm_scoreboard;
  `uvm_component_utils(apb_scoreboard)

  // Analysis implementation
  uvm_analysis_imp #(apb_seq_item, apb_scoreboard) analysis_imp;

  // Reference memory model
  bit [APB_DATA_W-1:0] ref_mem [256];

  // Statistics
  int unsigned checks_pass;
  int unsigned checks_fail;

  function new(string name = "apb_scoreboard", uvm_component parent = null);
    super.new(name, parent);
    analysis_imp = new("analysis_imp", this);
    checks_pass = 0;
    checks_fail = 0;
    // Initialize memory
    for (int i = 0; i < 256; i++) begin
      ref_mem[i] = 32'hDEADBEEF;
    end
  endfunction

  virtual function void write(apb_seq_item item);
    automatic int idx = item.addr[9:2];

    if (item.resp == APB_ERROR) begin
      `uvm_info("SCB", "Transaction with error response - not checking", UVM_MEDIUM)
      return;
    end

    if (item.dir == APB_WRITE) begin
      // Update reference model
      if (item.strb[0]) ref_mem[idx][7:0]   = item.wdata[7:0];
      if (item.strb[1]) ref_mem[idx][15:8]  = item.wdata[15:8];
      if (item.strb[2]) ref_mem[idx][23:16] = item.wdata[23:16];
      if (item.strb[3]) ref_mem[idx][31:24] = item.wdata[31:24];
      checks_pass++;
      `uvm_info("SCB", $sformatf("Write OK: %s", item.convert2string()), UVM_MEDIUM)
    end else begin
      // Check read data
      if (item.rdata == ref_mem[idx]) begin
        checks_pass++;
        `uvm_info("SCB", $sformatf("Read OK: %s", item.convert2string()), UVM_MEDIUM)
      end else begin
        checks_fail++;
        `uvm_error("SCB", $sformatf("Read MISMATCH: got=0x%08h exp=0x%08h",
                                    item.rdata, ref_mem[idx]))
      end
    end
  endfunction

  function void report_phase(uvm_phase phase);
    super.report_phase(phase);
    `uvm_info("SCB", $sformatf("Checks: %0d passed, %0d failed",
                               checks_pass, checks_fail), UVM_LOW)
    if (checks_fail == 0) begin
      `uvm_info("SCB", "*** TEST PASSED ***", UVM_NONE)
    end else begin
      `uvm_error("SCB", "*** TEST FAILED ***")
    end
  endfunction

endclass : apb_scoreboard

//===----------------------------------------------------------------------===//
// Environment: APB Verification Environment
//===----------------------------------------------------------------------===//

class apb_env extends uvm_env;
  `uvm_component_utils(apb_env)

  // Components
  apb_agent      agent;
  apb_scoreboard scoreboard;

  function new(string name = "apb_env", uvm_component parent = null);
    super.new(name, parent);
  endfunction

  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    agent      = apb_agent::type_id::create("agent", this);
    scoreboard = apb_scoreboard::type_id::create("scoreboard", this);
  endfunction

  virtual function void connect_phase(uvm_phase phase);
    super.connect_phase(phase);
    // Connect monitor to scoreboard
    agent.monitor.analysis_port.connect(scoreboard.analysis_imp);
  endfunction

endclass : apb_env

//===----------------------------------------------------------------------===//
// Test: APB Base Test
//===----------------------------------------------------------------------===//

class apb_base_test extends uvm_test;
  `uvm_component_utils(apb_base_test)

  apb_env env;

  function new(string name = "apb_base_test", uvm_component parent = null);
    super.new(name, parent);
  endfunction

  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    env = apb_env::type_id::create("env", this);
  endfunction

  virtual task run_phase(uvm_phase phase);
    apb_base_seq seq;

    phase.raise_objection(this);
    `uvm_info("TEST", "Starting APB base test", UVM_LOW)

    seq = apb_base_seq::type_id::create("seq");
    seq.num_txns = 10;
    seq.start(env.agent.sequencer);

    #100;
    `uvm_info("TEST", "APB base test complete", UVM_LOW)
    phase.drop_objection(this);
  endtask

  function void report_phase(uvm_phase phase);
    super.report_phase(phase);
    `uvm_info("TEST", "=== APB AVIP E2E Test Complete ===", UVM_NONE)
  endfunction

endclass : apb_base_test

//===----------------------------------------------------------------------===//
// Simple Memory DUT (for simulation)
//===----------------------------------------------------------------------===//

module apb_memory (
  input  logic                  clk,
  input  logic                  rst_n,
  input  logic [APB_ADDR_W-1:0] paddr,
  input  logic                  pselx,
  input  logic                  penable,
  input  logic                  pwrite,
  input  logic [APB_DATA_W-1:0] pwdata,
  input  logic [APB_STRB_W-1:0] pstrb,
  output logic [APB_DATA_W-1:0] prdata,
  output logic                  pready,
  output logic                  pslverr
);

  // Memory array
  logic [APB_DATA_W-1:0] mem [256];

  // Initialize memory
  initial begin
    for (int i = 0; i < 256; i++) begin
      mem[i] = 32'hDEADBEEF;
    end
  end

  // Always ready (no wait states)
  assign pready  = 1'b1;
  assign pslverr = 1'b0;

  // Memory read
  assign prdata = mem[paddr[9:2]];

  // Memory write
  always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
      // Reset handled by initial block
    end else if (pselx && penable && pwrite) begin
      if (pstrb[0]) mem[paddr[9:2]][7:0]   <= pwdata[7:0];
      if (pstrb[1]) mem[paddr[9:2]][15:8]  <= pwdata[15:8];
      if (pstrb[2]) mem[paddr[9:2]][23:16] <= pwdata[23:16];
      if (pstrb[3]) mem[paddr[9:2]][31:24] <= pwdata[31:24];
    end
  end

endmodule : apb_memory

//===----------------------------------------------------------------------===//
// Testbench Top Module
//===----------------------------------------------------------------------===//

module avip_e2e_tb;

  // Clock and reset
  logic clk;
  logic rst_n;

  // Clock generation
  initial begin
    clk = 0;
    forever #5 clk = ~clk;
  end

  // Reset generation
  initial begin
    rst_n = 0;
    #20 rst_n = 1;
  end

  // APB interface instance
  apb_if apb_bus (clk, rst_n);

  // DUT instance
  apb_memory dut (
    .clk     (clk),
    .rst_n   (rst_n),
    .paddr   (apb_bus.paddr),
    .pselx   (apb_bus.pselx),
    .penable (apb_bus.penable),
    .pwrite  (apb_bus.pwrite),
    .pwdata  (apb_bus.pwdata),
    .pstrb   (apb_bus.pstrb),
    .prdata  (apb_bus.prdata),
    .pready  (apb_bus.pready),
    .pslverr (apb_bus.pslverr)
  );

  // UVM test entry point
  initial begin
    // Set virtual interface in config_db (using full interface)
    uvm_config_db#(virtual apb_if)::set(null, "*", "vif", apb_bus);

    // Print test banner
    $display("========================================");
    $display("  AVIP E2E Testbench - Iteration 63");
    $display("========================================");

    // Run test
    run_test("apb_base_test");
  end

  // Timeout watchdog
  initial begin
    #10000;
    $display("ERROR: Test timeout!");
    $finish;
  end

endmodule : avip_e2e_tb

// PARSE: }
// MOORE: }

//===----------------------------------------------------------------------===//
// End of AVIP E2E Testbench
//===----------------------------------------------------------------------===//
