package alpha_pkg;
endpackage
