// RUN: circt-verilog --no-uvm-auto-include --ir-moore %s | FileCheck %s

module DPIOpenArraySupported;
  import "DPI-C" function void dpi_open_inout(
    input byte unsigned msg[],
    output byte unsigned digest[]
  );

  byte unsigned msg[];
  byte unsigned digest[];

  initial begin
    msg = new[2];
    msg[0] = 8'h12;
    msg[1] = 8'h34;
    digest = new[2];

    // Exercise call lowering with both input and output open-array arguments.
    dpi_open_inout(msg, digest);
    if (digest.size() != 2) begin
      $fatal(1, "unexpected digest size");
    end
  end

  // CHECK: %[[IN:.*]] = moore.read %msg : <open_uarray<i8>>
  // CHECK: %[[OUT_REF:.*]] = moore.variable : <open_uarray<i8>>
  // CHECK: func.call @dpi_open_inout(%[[IN]], %[[OUT_REF]]) : (!moore.open_uarray<i8>, !moore.ref<open_uarray<i8>>) -> ()
  // CHECK: %[[OUT_VAL:.*]] = moore.read %[[OUT_REF]] : <open_uarray<i8>>
  // CHECK: moore.blocking_assign %digest, %[[OUT_VAL]] : open_uarray<i8>
  // CHECK: func.func private @dpi_open_inout(!moore.open_uarray<i8>, !moore.ref<open_uarray<i8>>)
endmodule
