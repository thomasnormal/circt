`ifndef UVM_MACROS_SVH
`define UVM_MACROS_SVH
`endif
