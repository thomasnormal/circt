module always_ff;
endmodule
