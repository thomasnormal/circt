// RUN: circt-verilog --no-uvm-auto-include --ir-moore %s | FileCheck %s
// RUN: circt-verilog --no-uvm-auto-include --ir-moore %s

module SVABoundedAlwaysProperty(input logic clk, a, b, c, d);
  property p;
    @(posedge clk) a |-> b;
  endproperty

  // CHECK: %[[TRUE:.*]] = hw.constant true
  // CHECK: %[[D1:.*]] = ltl.delay %[[TRUE]], 1, 0 : i1
  // CHECK: %[[P1:.*]] = ltl.implication %[[D1]], %{{.*}} : !ltl.sequence, !ltl.property
  // CHECK: %[[D2:.*]] = ltl.delay %[[TRUE]], 2, 0 : i1
  // CHECK: %[[P2:.*]] = ltl.implication %[[D2]], %{{.*}} : !ltl.sequence, !ltl.property
  // CHECK: %[[AND1:.*]] = ltl.and %{{.*}}, %[[P1]], %[[P2]]
  // CHECK: verif.assert %[[AND1]] : !ltl.property
  assert property (always [0:2] p);

  // CHECK: %[[SPA:.*]] = ltl.and %[[D1]], %[[P1]] : !ltl.sequence, !ltl.property
  // CHECK: %[[SPB:.*]] = ltl.and %[[D2]], %[[P2]] : !ltl.sequence, !ltl.property
  // CHECK: %[[AND2:.*]] = ltl.and %[[SPA]], %[[SPB]] : !ltl.property, !ltl.property
  // CHECK: verif.assert %[[AND2]] : !ltl.property
  assert property (s_always [1:2] p);

  assert property (@(posedge clk) c |-> d);
endmodule
