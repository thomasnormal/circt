// RUN: circt-verilog %s --ir-hw -o %t.mlir
// RUN: circt-bmc --run-smtlib --ignore-asserts-until=1 -b 8 --module top %t.mlir | FileCheck %s

module top(input logic clk);
  logic [1:0] v = 2'b00;
  logic [2:0] step = 3'd0;

  always_ff @(posedge clk) begin
    case (step)
      3'd0: begin
        v <= 2'b10; // bit0 stays 0
        step <= 3'd1;
      end
      3'd1: begin
        v <= 2'b11; // bit0 rises 0->1
        step <= 3'd2;
      end
      3'd2: begin
        v <= 2'b01; // bit0 stays 1
        step <= 3'd3;
      end
      3'd3: begin
        v <= 2'b00; // bit0 falls 1->0
        step <= 3'd4;
      end
      3'd4: begin
        step <= 3'd5;
      end
      default: begin
        v <= v;
        step <= step;
      end
    endcase
  end

  assert property (@(posedge clk) (step == 3'd1) |-> !$rose(v));
  assert property (@(posedge clk) (step == 3'd2) |-> $rose(v));
  assert property (@(posedge clk) (step == 3'd3) |-> !$fell(v));
  assert property (@(posedge clk) (step == 3'd4) |-> $fell(v));
endmodule

// CHECK: BMC_RESULT=UNSAT
