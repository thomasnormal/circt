package uvm_pkg;
endpackage
