// Wrapper to ensure prim_ascon_duplex sees prim_flop_macros definitions.
`include "prim_flop_macros.sv"
`include "prim_ascon_duplex.sv"
