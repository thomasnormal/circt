module helper;
endmodule
