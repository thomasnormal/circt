module alpha;
endmodule

interface alpha_if;
endinterface

class alpha_cls;
endclass

program alpha_prog;
endprogram

checker alpha_chk;
endchecker
