// RUN: circt-verilog --ir-hw %s | \
// RUN:   circt-bmc --run-smtlib -b 4 --module=sva_concat_repeat_delay_range_unsat - | FileCheck %s
// REQUIRES: slang
// REQUIRES: z3

module sva_concat_repeat_delay_range_unsat(input logic clk);
  logic req;
  logic a;
  logic b;
  logic c;
  initial req = 1'b1;
  always @(posedge clk) begin
    req <= 1'b0;
  end
  assign a = 1'b1;
  assign b = 1'b1;
  assign c = 1'b1;
  assert property (@(posedge clk) req |-> (a ##1 b) [*2] ##[1:2] c);
endmodule

// CHECK: BMC_RESULT=UNSAT
