`include "legacy.sv"
module top;
endmodule
