// Wrapper to inject prim_assert macros for usb_fs_tx.
`include "prim_assert.sv"
`include "usb_fs_tx.sv"
