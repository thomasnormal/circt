// Wrapper to inject prim_assert macros for usbdev_linkstate.
`include "prim_assert.sv"
`include "usbdev_linkstate.sv"
