package SpiMasterPkg;
  `include "SpiMasterSeqItemConverter.sv"
endpackage
