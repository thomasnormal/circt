// Wrapper to inject prim_assert macros for spi_host_fsm.
`include "prim_assert.sv"
`include "spi_host_fsm.sv"
