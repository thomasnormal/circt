// Wrapper to inject prim_assert macros for usbdev_usbif.
`include "prim_assert.sv"
`include "usbdev_usbif.sv"
