`ifdef HELLO
import hello::defined;
`else
import hello::undefined;
`endif
