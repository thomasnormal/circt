package DummyReadEnvPkg;
endpackage
