`define WHICH include_cfg_mod
