package DummySlaveReadEnvPkg;
endpackage
